package jtag;

typedef enum logic [3:0] {
    TEST_LOGIC_RESET, RUN_TEST_IDLE, SELECT_DR_SCAN, CAPTURE_DR, SHIFT_DR,
    EXIT1_DR, PAUSE_DR, EXIT2_DR, UPDATE_DR, SELECT_IR_SCAN, CAPTURE_IR,
    SHIFT_IR, EXIT1_IR, PAUSE_IR, EXIT2_IR, UPDATE_IR
} jtag_state_t;

endpackage