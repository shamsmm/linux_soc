//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Thu Jun  5 19:29:35 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [31:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire [15:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b1;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0008000180002000C0000E002300020062002000620200006200000802000030;
defparam prom_inst_0.INIT_RAM_01 = 256'h000000000000000000000000DFFB0EFEFEFF0500620000000EFEFEFF05006200;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[15:0],dout[31:16]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b1;
defparam prom_inst_1.BIT_WIDTH = 16;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h130313056F0013056F00630413FE83A323A8130323AC130323A613039382B702;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000000000000000000006FF0E39E938E930E23A41303E39E938E930E23A4;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_pROM
